`timescale 1ns/1ps

module breathing_water_led (
    input  wire        clk,              
    input  wire        rst,              
    input  wire        dip_switch_mode,  
    output reg [15:0]  led               
);

    // === �������� ===
    localparam CLK_FREQ        = 100_000_000;    // 100MHz
    localparam PWM_FREQ        = 1000;           // 1KHz PWM
    localparam PWM_PERIOD      = CLK_FREQ / PWM_FREQ;           // 100_000
    localparam BREATH_STEP_CNT = 100;            // ����100��
    localparam BREATH_TOTAL_MS = 8000;           // ����8������
    localparam BREATH_CNT_STEP = BREATH_TOTAL_MS / (BREATH_STEP_CNT*2); // 8s/200��
    localparam BREATH_STEP_CLK = (CLK_FREQ/1000) * BREATH_CNT_STEP; // ÿ������ʱ��

    // === ״̬�Ĵ������� ===
    reg [$clog2(PWM_PERIOD)-1:0]     pwm_cnt = 0;               // PWM����
    reg [$clog2(BREATH_STEP_CLK)-1:0] breath_time_cnt = 0;      // ����step����
    reg [6:0]                        breath_step = 0;           // ��ǰ���ȵȼ�
    reg                              breath_up = 1;             // ��������

    // ---- ��ˮ������ר��
    reg [3:0]   led_main = 0;      // ��ǰ����LED
    reg [3:0]   led_fade = 0;      // ��һ������LED
    reg [6:0]   bright_main = 0;   // ���ڱ���LED����
    reg [6:0]   bright_fade = 0;   // ����LED����
    reg         fw_dir = 0;        // ��������0��/1��
    reg [31:0]  water_timer = 0;   // ������ʱ

    // === ���뿪�ؿ���ģʽ ===
    wire fn_mode = dip_switch_mode; // ������ƹ����л���0Ϊ�����ƣ�1Ϊ��ˮ��

    // === ���������ȣ�����1�� ===
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            breath_step     <= 0;
            breath_up       <= 1;
            breath_time_cnt <= 0;
        end else if (!fn_mode) begin
            // ���ں�����ģʽ�¹���
            if (breath_time_cnt < BREATH_STEP_CLK - 1)
                breath_time_cnt <= breath_time_cnt + 1;
            else begin
                breath_time_cnt <= 0;
                if (breath_up) begin
                    if (breath_step < BREATH_STEP_CNT)
                        breath_step <= breath_step + 1;
                    else
                        breath_up <= 0;
                end else begin
                    if (breath_step > 0)
                        breath_step <= breath_step - 1;
                    else
                        breath_up <= 1;
                end
            end
        end
    end

    // === PWM������ ===
    always @(posedge clk or posedge rst) begin
        if (rst)
            pwm_cnt <= 0;
        else if (pwm_cnt < PWM_PERIOD - 1)
            pwm_cnt <= pwm_cnt + 1;
        else
            pwm_cnt <= 0;
    end

    // === ��ˮ�����߼�������2�� ===
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            led_main    <= 0;
            led_fade    <= 0;
            bright_main <= 0;
            bright_fade <= 0;
            fw_dir      <= 0;
            water_timer <= 0;
        end else if (fn_mode) begin
            if (water_timer < BREATH_STEP_CLK-1)
                water_timer <= water_timer + 1;
            else begin
                water_timer <= 0;
                // ��LED����
                if (bright_main < BREATH_STEP_CNT)
                    bright_main <= bright_main + 1;
                // ����LED�䰵
                if (bright_fade > 0)
                    bright_fade <= bright_fade - 1;

                // ��LED������������һλ������һλfade
                if (bright_main == BREATH_STEP_CNT) begin
                    led_fade     <= led_main;        // ��ǰλתΪ����
                    bright_fade  <= BREATH_STEP_CNT; // ������������
                    // �ı���LEDλ��
                    if (!fw_dir) begin
                        if (led_main < 15)
                            led_main <= led_main + 1;
                        else begin
                            led_main <= 14;
                            fw_dir   <= 1;
                        end
                    end else begin
                        if (led_main > 0)
                            led_main <= led_main - 1;
                        else begin
                            led_main <= 1;
                            fw_dir <= 0;
                        end
                    end
                    bright_main <= 0; // ����LED��0��ʼ����
                end
            end
        end
    end

    // === PWM������� ===
    reg [15:0] led_pwm;
    always @(posedge clk or posedge rst) begin
        if (rst)
            led <= 16'b0;
        else if (!fn_mode) begin
            // ����1��������ģʽ����8����8����
            // ��8������������8�����½�
            if (pwm_cnt < breath_step * PWM_PERIOD / BREATH_STEP_CNT)
                led[7:0] <= 8'hFF;
            else
                led[7:0] <= 8'h00;
            if (pwm_cnt < (BREATH_STEP_CNT-breath_step) * PWM_PERIOD / BREATH_STEP_CNT)
                led[15:8] <= 8'hFF;
            else
                led[15:8] <= 8'h00;
        end else begin
            // ����2����ˮ����ģʽ���������Ƚ����ص�
            led_pwm = 16'b0;
            if (pwm_cnt < (bright_main * PWM_PERIOD / BREATH_STEP_CNT))
                led_pwm[led_main] = 1'b1;
            if (bright_fade > 0 && (led_fade != led_main))
                if (pwm_cnt < (bright_fade * PWM_PERIOD / BREATH_STEP_CNT))
                    led_pwm[led_fade] = 1'b1;
            led <= led_pwm;
        end
    end

endmodule
